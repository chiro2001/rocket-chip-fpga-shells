// name cc_dir_ext depth 256 width 34 ports mrw mask_gran 17 
// name cc_banks_0_ext depth 4096 width 32 ports rw  
// name data_arrays_0_ext depth 4096 width 32 ports mrw mask_gran 8 
// name tag_array_ext depth 256 width 20 ports rw  
// name tag_array_0_ext depth 256 width 19 ports mrw mask_gran 19 
// name data_arrays_0_0_ext depth 4096 width 32 ports mrw mask_gran 32 

`define DRM \
  .wr_data(RW0_wdata),\
  .wr_addr(RW0_addr),\
  .wr_en(RW0_wmode & RW0_en & RW0_wmask),\
  .wr_clk(RW0_clk),\
  .wr_rst(0),\
  .rd_addr(RW0_addr),\
  .rd_data(RW0_rdata),\
  .rd_clk(rd_clk),\
  .rd_rst(0)

`define DRMM \
  .wr_data(RW0_wdata),\
  .wr_addr(RW0_addr),\
  .wr_en(RW0_wmode & RW0_en),\
  .wr_byte_en(RW0_wmask),\
  .wr_clk(RW0_clk),\
  .wr_rst(0),\
  .rd_addr(RW0_addr),\
  .rd_data(RW0_rdata),\
  .rd_clk(rd_clk),\
  .rd_rst(0)

module split_drm_36x128(
  input  [6:0]  RW0_addr,
  input         RW0_clk,
  input  [31:0] RW0_wdata,
  output [31:0] RW0_rdata,
  input         RW0_en,
  input         RW0_wmode,
  input         RW0_wmask
);
drm_36x128 inst (`DRMM);
endmodule

module split_drm_8x1024(
  input  [9:0]  RW0_addr,
  input         RW0_clk,
  input  [7:0]  RW0_wdata,
  output [7:0]  RW0_rdata,
  input         RW0_en,
  input         RW0_wmode,
  input         RW0_wmask
);
drm_8x1024 drm_8x1024_inst (`DRMM);
endmodule

module split_drm_15x1024(
  input  [9:0]  RW0_addr,
  input         RW0_clk,
  input  [14:0] RW0_wdata,
  output [14:0] RW0_rdata,
  input         RW0_en,
  input         RW0_wmode,
  input         RW0_wmask
);
wire [7:0] RW0_rdata_0;
wire [6:0] RW0_rdata_1;
assign RW0_rdata = {RW0_rdata_1, RW0_rdata_0};
split_drm_8x1024 split_drm_8x1024_inst_0 (
  .RW0_addr(RW0_addr),
  .RW0_clk(RW0_clk),
  .RW0_wdata(RW0_wdata[7:0]),
  .RW0_rdata(RW0_rdata_0),
  .RW0_en(RW0_en),
  .RW0_wmode(RW0_wmode),
  .RW0_wmask(RW0_wmask)
);
split_drm_8x1024 split_drm_8x1024_inst_1 (
  .RW0_addr(RW0_addr),
  .RW0_clk(RW0_clk),
  .RW0_wdata(RW0_wdata[14:8]),
  .RW0_rdata(RW0_rdata_1),
  .RW0_en(RW0_en),
  .RW0_wmode(RW0_wmode),
  .RW0_wmask(RW0_wmask)
);
endmodule

module split_drm_32x1024_nomask(
  input  [9:0]    RW0_addr,
  input           RW0_clk,
  input  [31:0]   RW0_wdata,
  output [31:0]   RW0_rdata,
  input           RW0_en,
  input           RW0_wmode,
  input           RW0_wmask
);
drm_32x1024 inst (`DRM);
endmodule

module split_drm_32x1024(
  input  [9:0]    RW0_addr,
  input           RW0_clk,
  input  [31:0]   RW0_wdata,
  output [31:0]   RW0_rdata,
  input           RW0_en,
  input           RW0_wmode,
  input  [7:0]    RW0_wmask
);
  wire [11:0] mem_0_0_RW0_addr;
  wire  mem_0_0_RW0_clk;
  wire [7:0] mem_0_0_RW0_wdata;
  wire [7:0] mem_0_0_RW0_rdata;
  wire  mem_0_0_RW0_en;
  wire  mem_0_0_RW0_wmode;
  wire  mem_0_0_RW0_wmask;
  wire [11:0] mem_0_1_RW0_addr;
  wire  mem_0_1_RW0_clk;
  wire [7:0] mem_0_1_RW0_wdata;
  wire [7:0] mem_0_1_RW0_rdata;
  wire  mem_0_1_RW0_en;
  wire  mem_0_1_RW0_wmode;
  wire  mem_0_1_RW0_wmask;
  wire [11:0] mem_0_2_RW0_addr;
  wire  mem_0_2_RW0_clk;
  wire [7:0] mem_0_2_RW0_wdata;
  wire [7:0] mem_0_2_RW0_rdata;
  wire  mem_0_2_RW0_en;
  wire  mem_0_2_RW0_wmode;
  wire  mem_0_2_RW0_wmask;
  wire [11:0] mem_0_3_RW0_addr;
  wire  mem_0_3_RW0_clk;
  wire [7:0] mem_0_3_RW0_wdata;
  wire [7:0] mem_0_3_RW0_rdata;
  wire  mem_0_3_RW0_en;
  wire  mem_0_3_RW0_wmode;
  wire  mem_0_3_RW0_wmask;
  wire [7:0] RW0_rdata_0_0 = mem_0_0_RW0_rdata;
  wire [7:0] RW0_rdata_0_1 = mem_0_1_RW0_rdata;
  wire [7:0] RW0_rdata_0_2 = mem_0_2_RW0_rdata;
  wire [7:0] RW0_rdata_0_3 = mem_0_3_RW0_rdata;
  wire [15:0] _GEN_0 = {RW0_rdata_0_1,RW0_rdata_0_0};
  wire [23:0] _GEN_1 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [31:0] RW0_rdata_0 = {RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [15:0] _GEN_2 = {RW0_rdata_0_1,RW0_rdata_0_0};
  wire [23:0] _GEN_3 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  split_drm_8x1024 mem_0_0 (
    .RW0_addr(mem_0_0_RW0_addr),
    .RW0_clk(mem_0_0_RW0_clk),
    .RW0_wdata(mem_0_0_RW0_wdata),
    .RW0_rdata(mem_0_0_RW0_rdata),
    .RW0_en(mem_0_0_RW0_en),
    .RW0_wmode(mem_0_0_RW0_wmode),
    .RW0_wmask(mem_0_0_RW0_wmask)
  );
  split_drm_8x1024 mem_0_1 (
    .RW0_addr(mem_0_1_RW0_addr),
    .RW0_clk(mem_0_1_RW0_clk),
    .RW0_wdata(mem_0_1_RW0_wdata),
    .RW0_rdata(mem_0_1_RW0_rdata),
    .RW0_en(mem_0_1_RW0_en),
    .RW0_wmode(mem_0_1_RW0_wmode),
    .RW0_wmask(mem_0_1_RW0_wmask)
  );
  split_drm_8x1024 mem_0_2 (
    .RW0_addr(mem_0_2_RW0_addr),
    .RW0_clk(mem_0_2_RW0_clk),
    .RW0_wdata(mem_0_2_RW0_wdata),
    .RW0_rdata(mem_0_2_RW0_rdata),
    .RW0_en(mem_0_2_RW0_en),
    .RW0_wmode(mem_0_2_RW0_wmode),
    .RW0_wmask(mem_0_2_RW0_wmask)
  );
  split_drm_8x1024 mem_0_3 (
    .RW0_addr(mem_0_3_RW0_addr),
    .RW0_clk(mem_0_3_RW0_clk),
    .RW0_wdata(mem_0_3_RW0_wdata),
    .RW0_rdata(mem_0_3_RW0_rdata),
    .RW0_en(mem_0_3_RW0_en),
    .RW0_wmode(mem_0_3_RW0_wmode),
    .RW0_wmask(mem_0_3_RW0_wmask)
  );
  assign RW0_rdata = {RW0_rdata_0_3,_GEN_1};
  assign mem_0_0_RW0_addr = RW0_addr;
  assign mem_0_0_RW0_clk = RW0_clk;
  assign mem_0_0_RW0_wdata = RW0_wdata[7:0];
  assign mem_0_0_RW0_en = RW0_en;
  assign mem_0_0_RW0_wmode = RW0_wmode;
  assign mem_0_0_RW0_wmask = RW0_wmask;
  assign mem_0_1_RW0_addr = RW0_addr;
  assign mem_0_1_RW0_clk = RW0_clk;
  assign mem_0_1_RW0_wdata = RW0_wdata[15:8];
  assign mem_0_1_RW0_en = RW0_en;
  assign mem_0_1_RW0_wmode = RW0_wmode;
  assign mem_0_1_RW0_wmask = RW0_wmask;
  assign mem_0_2_RW0_addr = RW0_addr;
  assign mem_0_2_RW0_clk = RW0_clk;
  assign mem_0_2_RW0_wdata = RW0_wdata[23:16];
  assign mem_0_2_RW0_en = RW0_en;
  assign mem_0_2_RW0_wmode = RW0_wmode;
  assign mem_0_2_RW0_wmask = RW0_wmask;
  assign mem_0_3_RW0_addr = RW0_addr;
  assign mem_0_3_RW0_clk = RW0_clk;
  assign mem_0_3_RW0_wdata = RW0_wdata[31:24];
  assign mem_0_3_RW0_en = RW0_en;
  assign mem_0_3_RW0_wmode = RW0_wmode;
  assign mem_0_3_RW0_wmask = RW0_wmask;
endmodule

module split_drm_128x1024(
  input  [9:0]    RW0_addr,
  input           RW0_clk,
  input  [127:0]  RW0_wdata,
  output [127:0]  RW0_rdata,
  input           RW0_en,
  input           RW0_wmode,
  input           RW0_wmask
);
  wire [11:0] mem_0_0_RW0_addr;
  wire  mem_0_0_RW0_clk;
  wire [31:0] mem_0_0_RW0_wdata;
  wire [31:0] mem_0_0_RW0_rdata;
  wire  mem_0_0_RW0_en;
  wire  mem_0_0_RW0_wmode;
  wire  mem_0_0_RW0_wmask;
  wire [11:0] mem_0_1_RW0_addr;
  wire  mem_0_1_RW0_clk;
  wire [31:0] mem_0_1_RW0_wdata;
  wire [31:0] mem_0_1_RW0_rdata;
  wire  mem_0_1_RW0_en;
  wire  mem_0_1_RW0_wmode;
  wire  mem_0_1_RW0_wmask;
  wire [11:0] mem_0_2_RW0_addr;
  wire  mem_0_2_RW0_clk;
  wire [31:0] mem_0_2_RW0_wdata;
  wire [31:0] mem_0_2_RW0_rdata;
  wire  mem_0_2_RW0_en;
  wire  mem_0_2_RW0_wmode;
  wire  mem_0_2_RW0_wmask;
  wire [11:0] mem_0_3_RW0_addr;
  wire  mem_0_3_RW0_clk;
  wire [31:0] mem_0_3_RW0_wdata;
  wire [31:0] mem_0_3_RW0_rdata;
  wire  mem_0_3_RW0_en;
  wire  mem_0_3_RW0_wmode;
  wire  mem_0_3_RW0_wmask;
  wire [31:0] RW0_rdata_0_0 = mem_0_0_RW0_rdata;
  wire [31:0] RW0_rdata_0_1 = mem_0_1_RW0_rdata;
  wire [31:0] RW0_rdata_0_2 = mem_0_2_RW0_rdata;
  wire [31:0] RW0_rdata_0_3 = mem_0_3_RW0_rdata;
  wire [15:0] _GEN_0 = {RW0_rdata_0_1,RW0_rdata_0_0};
  wire [23:0] _GEN_1 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [31:0] RW0_rdata_0 = {RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [15:0] _GEN_2 = {RW0_rdata_0_1,RW0_rdata_0_0};
  wire [23:0] _GEN_3 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  split_drm_32x1024 mem_0_0 (
    .RW0_addr(mem_0_0_RW0_addr),
    .RW0_clk(mem_0_0_RW0_clk),
    .RW0_wdata(mem_0_0_RW0_wdata),
    .RW0_rdata(mem_0_0_RW0_rdata),
    .RW0_en(mem_0_0_RW0_en),
    .RW0_wmode(mem_0_0_RW0_wmode),
    .RW0_wmask(mem_0_0_RW0_wmask)
  );
  split_drm_32x1024 mem_0_1 (
    .RW0_addr(mem_0_1_RW0_addr),
    .RW0_clk(mem_0_1_RW0_clk),
    .RW0_wdata(mem_0_1_RW0_wdata),
    .RW0_rdata(mem_0_1_RW0_rdata),
    .RW0_en(mem_0_1_RW0_en),
    .RW0_wmode(mem_0_1_RW0_wmode),
    .RW0_wmask(mem_0_1_RW0_wmask)
  );
  split_drm_32x1024 mem_0_2 (
    .RW0_addr(mem_0_2_RW0_addr),
    .RW0_clk(mem_0_2_RW0_clk),
    .RW0_wdata(mem_0_2_RW0_wdata),
    .RW0_rdata(mem_0_2_RW0_rdata),
    .RW0_en(mem_0_2_RW0_en),
    .RW0_wmode(mem_0_2_RW0_wmode),
    .RW0_wmask(mem_0_2_RW0_wmask)
  );
  split_drm_32x1024 mem_0_3 (
    .RW0_addr(mem_0_3_RW0_addr),
    .RW0_clk(mem_0_3_RW0_clk),
    .RW0_wdata(mem_0_3_RW0_wdata),
    .RW0_rdata(mem_0_3_RW0_rdata),
    .RW0_en(mem_0_3_RW0_en),
    .RW0_wmode(mem_0_3_RW0_wmode),
    .RW0_wmask(mem_0_3_RW0_wmask)
  );
  assign RW0_rdata = {RW0_rdata_0_3,_GEN_1};
  assign mem_0_0_RW0_addr = RW0_addr;
  assign mem_0_0_RW0_clk = RW0_clk;
  assign mem_0_0_RW0_wdata = RW0_wdata[31:0];
  assign mem_0_0_RW0_en = RW0_en;
  assign mem_0_0_RW0_wmode = RW0_wmode;
  assign mem_0_0_RW0_wmask = RW0_wmask;
  assign mem_0_1_RW0_addr = RW0_addr;
  assign mem_0_1_RW0_clk = RW0_clk;
  assign mem_0_1_RW0_wdata = RW0_wdata[63:32];
  assign mem_0_1_RW0_en = RW0_en;
  assign mem_0_1_RW0_wmode = RW0_wmode;
  assign mem_0_1_RW0_wmask = RW0_wmask;
  assign mem_0_2_RW0_addr = RW0_addr;
  assign mem_0_2_RW0_clk = RW0_clk;
  assign mem_0_2_RW0_wdata = RW0_wdata[95:64];
  assign mem_0_2_RW0_en = RW0_en;
  assign mem_0_2_RW0_wmode = RW0_wmode;
  assign mem_0_2_RW0_wmask = RW0_wmask;
  assign mem_0_3_RW0_addr = RW0_addr;
  assign mem_0_3_RW0_clk = RW0_clk;
  assign mem_0_3_RW0_wdata = RW0_wdata[127:96];
  assign mem_0_3_RW0_en = RW0_en;
  assign mem_0_3_RW0_wmode = RW0_wmode;
  assign mem_0_3_RW0_wmask = RW0_wmask;
endmodule

module split_drm_17x256(
  input  [7:0]    RW0_addr,
  input           RW0_clk,
  input  [16:0]   RW0_wdata,
  output [16:0]   RW0_rdata,
  input           RW0_en,
  input           RW0_wmode,
  input           RW0_wmask
);
drm_17x256 inst (`DRM);
endmodule
module split_drm_32x4096(
  input  [11:0]   RW0_addr,
  input           RW0_clk,
  input  [31:0]   RW0_wdata,
  output [31:0]   RW0_rdata,
  input           RW0_en,
  input           RW0_wmode,
  input           RW0_wmask
);
drm_32x4096 inst (`DRM);
endmodule
module split_drm_8x4096(
  input  [11:0]   RW0_addr,
  input           RW0_clk,
  input  [7:0]    RW0_wdata,
  output [7:0]    RW0_rdata,
  input           RW0_en,
  input           RW0_wmode,
  input           RW0_wmask
);
drm_8x4096 inst (`DRM);
endmodule
module split_drm_20x256(
  input  [7:0]    RW0_addr,
  input           RW0_clk,
  input  [19:0]   RW0_wdata,
  output [19:0]   RW0_rdata,
  input           RW0_en,
  input           RW0_wmode,
  input           RW0_wmask
);
drm_20x256 inst (`DRM);
endmodule
module split_drm_21x64(
  input  [5:0]    RW0_addr,
  input           RW0_clk,
  input  [20:0]   RW0_wdata,
  output [20:0]   RW0_rdata,
  input           RW0_en,
  input           RW0_wmode,
  input           RW0_wmask
);
drm_21x64 inst (`DRM);
endmodule
module split_drm_64x8192(
  input  [12:0]   RW0_addr,
  input           RW0_clk,
  input  [63:0]   RW0_wdata,
  output [63:0]   RW0_rdata,
  input           RW0_en,
  input           RW0_wmode,
  input  [7:0]    RW0_wmask
);
drm_64x8192 inst (`DRMM);
endmodule
