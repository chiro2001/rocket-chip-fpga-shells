module split_data_arrays_0_ext(input [9:0] RW0_addr,
                               input RW0_clk,
                               input [7:0] RW0_wdata,
                               output [7:0] RW0_rdata,
                               input RW0_en,
                               input RW0_wmode,
                               input RW0_wmask);
wire wen;
assign wen = RW0_en & RW0_en & RW0_wmask;
GTP_DRM9K
#(
.DATA_WIDTH_A (8), // 1 2 4 8 16 32 9 18 36
.DATA_WIDTH_B (8), // 1 2 4 8 16 32 9 18 36
.WRITE_MODE_A ("NORMAL_WRITE"), // TRANSPARENT_WRITE READ_BEFORE_WRITE
.WRITE_MODE_B ("NORMAL_WRITE"), // TRANSPARENT_WRITE READ_BEFORE_WRITE
.DOA_REG (0),
.DOB_REG (0),
.RST_TYPE ("SYNC"), // ASYNC,ASYNC_SYNC_RELEASE
.RAM_MODE ("TRUE_DUAL_PORT"), // SIMPLE_DUAL_PORT SINGLE_PORT ROM
.GRS_EN ("TRUE"), //"TRUE"; "FALSE" 使能内部复位
.DOA_REG_CLKINV (1'b0), //clka polarity invert for output register
.DOB_REG_CLKINV (1'b0), //clkb polarity invert for output register
.INIT_00 (288'h000000000000000000000000000000000000000000000000000000000000000000000000),
.INIT_01 (288'h000000000000000000000000000000000000000000000000000000000000000000000000),
.INIT_02 (288'h000000000000000000000000000000000000000000000000000000000000000000000000),
.INIT_03 (288'h000000000000000000000000000000000000000000000000000000000000000000000000),
.INIT_04 (288'h000000000000000000000000000000000000000000000000000000000000000000000000),
.INIT_05 (288'h000000000000000000000000000000000000000000000000000000000000000000000000),
.INIT_06 (288'h000000000000000000000000000000000000000000000000000000000000000000000000),
.INIT_07 (288'h000000000000000000000000000000000000000000000000000000000000000000000000),
.INIT_08 (288'h000000000000000000000000000000000000000000000000000000000000000000000000),
.INIT_09 (288'h000000000000000000000000000000000000000000000000000000000000000000000000),
.INIT_0A (288'h000000000000000000000000000000000000000000000000000000000000000000000000),
.INIT_0B (288'h000000000000000000000000000000000000000000000000000000000000000000000000),
.INIT_0C (288'h000000000000000000000000000000000000000000000000000000000000000000000000),
.INIT_0D (288'h000000000000000000000000000000000000000000000000000000000000000000000000),
.INIT_0E (288'h000000000000000000000000000000000000000000000000000000000000000000000000),
.INIT_0F (288'h000000000000000000000000000000000000000000000000000000000000000000000000),
.INIT_10 (288'h000000000000000000000000000000000000000000000000000000000000000000000000),
.INIT_11 (288'h000000000000000000000000000000000000000000000000000000000000000000000000),
.INIT_12 (288'h000000000000000000000000000000000000000000000000000000000000000000000000),
.INIT_13 (288'h000000000000000000000000000000000000000000000000000000000000000000000000),
.INIT_14 (288'h000000000000000000000000000000000000000000000000000000000000000000000000),
.INIT_15 (288'h000000000000000000000000000000000000000000000000000000000000000000000000),
.INIT_16 (288'h000000000000000000000000000000000000000000000000000000000000000000000000),
.INIT_17 (288'h000000000000000000000000000000000000000000000000000000000000000000000000),
.INIT_18 (288'h000000000000000000000000000000000000000000000000000000000000000000000000),
.INIT_19 (288'h000000000000000000000000000000000000000000000000000000000000000000000000),
.INIT_1A (288'h000000000000000000000000000000000000000000000000000000000000000000000000),
.INIT_1B (288'h000000000000000000000000000000000000000000000000000000000000000000000000),
.INIT_1C (288'h000000000000000000000000000000000000000000000000000000000000000000000000),
.INIT_1D (288'h000000000000000000000000000000000000000000000000000000000000000000000000),
.INIT_1E (288'h000000000000000000000000000000000000000000000000000000000000000000000000),
.INIT_1F (288'h000000000000000000000000000000000000000000000000000000000000000000000000),
.INIT_FILE ("NONE"),
.SIM_DEVICE ("PGL22G")
//add for initialization memory
// .BLOCK_X (0) , //indicate X location of block memory when cascaded with DRM18Ks
// .BLOCK_Y (0) , //indicate Y location of block memory when cascaded with DRM18Ks
// .RAM_DATA_WIDTH (8), //the total DATA WIDTH of cascaded DRMS
// .RAM_ADDR_WIDTH (10), //the total ADDR WIDTH of cascaded DRMS
// .INIT_FORMAT ("BIN") //initial file data type binary or hexadecimal
)
// SDP RAM
GTP_DRM9K_inst (
/**
 WADDR ADDRA 输入 写地址输入
 DI DIA 输入 数据输入
 WE WEA 输入 写使能
 WCLK CLKA 输入 写时钟
 WCE CEA 输入 写时钟使能
 WRST RSTA 输入 写寄存器复位
 Q DOB 输出 数据输出
 RADDR ADDRB 输入 读地址输入
 RCLK CLKB 输入 读时钟
 RCE CEB 输入 读时钟使能
 RORCE ORCEB 输入 读出寄存器OE
 RRST RSTB 输入 读寄存器复位
 */
// .DOA (DOA),
.ADDRA (RW0_addr),
// .ADDRA_HOLD (ADDRA_HOLD),
.DIA (RW0_wdata),
.WEA (wen),
.CLKA (RW0_clk),
.CEA (1),
// .ORCEA (ORCEA),
// .RSTA (0),
.DOB (RW0_rdata),
.ADDRB (RW0_addr),
// .ADDRB_HOLD (ADDRB_HOLD),
// .DIB (DIB),
// .WEB (WEB),
.CLKB (RW0_clk),
.CEB (1),
// .ORCEB (ORCEB),
.ORCEB (0)
// .RSTB (RSTB)
);
endmodule
